`timescale  1ns / 1ns
// 1024x24 synchronous ROM with fixed (random) content
//
module  rom1024x24  (
  input  logic            clk ,  // Rising-edge clock
  input  logic            cen ,  // Chip-enable
  input  logic    [9:0]   adr ,  // Address input
  output logic    [23:0]  dout   // Data output
) ;

// Define ROM contents using case statement
//
always_ff  @ ( posedge clk )
  if  ( cen )
    case  ( adr )
		10'h0: dout <= #1 24'hFFF940;
		10'h1: dout <= #1 24'hAD0;
		10'h2: dout <= #1 24'hCCB;
		10'h3: dout <= #1 24'hFFFB55;
		10'h4: dout <= #1 24'hFFFAB1;
		10'h5: dout <= #1 24'hED;
		10'h6: dout <= #1 24'hF44;
		10'h7: dout <= #1 24'hA88;
		10'h8: dout <= #1 24'h8CD;
		10'h9: dout <= #1 24'h274;
		10'hA: dout <= #1 24'hFFF9F3;
		10'hB: dout <= #1 24'hD82;
		10'hC: dout <= #1 24'h3F9;
		10'hD: dout <= #1 24'hDEE;
		10'hE: dout <= #1 24'hFFF494;
		10'hF: dout <= #1 24'hFFF83B;
		10'h10: dout <= #1 24'h404;
		10'h11: dout <= #1 24'hFFF4E8;
		10'h12: dout <= #1 24'h308;
		10'h13: dout <= #1 24'hFFFF82;
		10'h14: dout <= #1 24'hFFF63E;
		10'h15: dout <= #1 24'hFFFF73;
		10'h16: dout <= #1 24'hFFFE1A;
		10'h17: dout <= #1 24'h359;
		10'h18: dout <= #1 24'h6D0;
		10'h19: dout <= #1 24'h39E;
		10'h1A: dout <= #1 24'hFFFD3D;
		10'h1B: dout <= #1 24'hFFFD27;
		10'h1C: dout <= #1 24'hFFFEF5;
		10'h1D: dout <= #1 24'h33;
		10'h1E: dout <= #1 24'hFFFA40;
		10'h1F: dout <= #1 24'hFFF566;
		10'h20: dout <= #1 24'hFFFAB4;
		10'h21: dout <= #1 24'hFFF15C;
		10'h22: dout <= #1 24'h861;
		10'h23: dout <= #1 24'hFFEE65;
		10'h24: dout <= #1 24'hFFF9A1;
		10'h25: dout <= #1 24'h3A7;
		10'h26: dout <= #1 24'h53A;
		10'h27: dout <= #1 24'h6F0;
		10'h28: dout <= #1 24'hFFF743;
		10'h29: dout <= #1 24'h20;
		10'h2A: dout <= #1 24'hFFF587;
		10'h2B: dout <= #1 24'hC2B;
		10'h2C: dout <= #1 24'h90B;
		10'h2D: dout <= #1 24'hFFFD1E;
		10'h2E: dout <= #1 24'h18B;
		10'h2F: dout <= #1 24'h275;
		10'h30: dout <= #1 24'hFFFA50;
		10'h31: dout <= #1 24'hFFFF44;
		10'h32: dout <= #1 24'hFFFAEA;
		10'h33: dout <= #1 24'h218;
		10'h34: dout <= #1 24'h264;
		10'h35: dout <= #1 24'h818;
		10'h36: dout <= #1 24'hFFF07A;
		10'h37: dout <= #1 24'h329;
		10'h38: dout <= #1 24'h353;
		10'h39: dout <= #1 24'hBA5;
		10'h3A: dout <= #1 24'hFFEB54;
		10'h3B: dout <= #1 24'hFFF358;
		10'h3C: dout <= #1 24'hFFFDF5;
		10'h3D: dout <= #1 24'h441;
		10'h3E: dout <= #1 24'hFFF5E3;
		10'h3F: dout <= #1 24'hFFF7C7;
		10'h40: dout <= #1 24'hFFFE2B;
		10'h41: dout <= #1 24'h3E2;
		10'h42: dout <= #1 24'hFFFC73;
		10'h43: dout <= #1 24'hD9;
		10'h44: dout <= #1 24'hFFFA40;
		10'h45: dout <= #1 24'h5D;
		10'h46: dout <= #1 24'hFFF52B;
		10'h47: dout <= #1 24'h4AB;
		10'h48: dout <= #1 24'h12E2;
		10'h49: dout <= #1 24'h722;
		10'h4A: dout <= #1 24'hFFF788;
		10'h4B: dout <= #1 24'hFFFCAA;
		10'h4C: dout <= #1 24'hFFF786;
		10'h4D: dout <= #1 24'hFFF4BC;
		10'h4E: dout <= #1 24'hFFEFCF;
		10'h4F: dout <= #1 24'h4EA;
		10'h50: dout <= #1 24'hFFF82F;
		10'h51: dout <= #1 24'hFFFEC6;
		10'h52: dout <= #1 24'hFFF5F2;
		10'h53: dout <= #1 24'hFFF6E2;
		10'h54: dout <= #1 24'hFFF9E0;
		10'h55: dout <= #1 24'hFFF8C9;
		10'h56: dout <= #1 24'hFFF9C9;
		10'h57: dout <= #1 24'hA01;
		10'h58: dout <= #1 24'hFFF9DD;
		10'h59: dout <= #1 24'h3C0;
		10'h5A: dout <= #1 24'h515;
		10'h5B: dout <= #1 24'hFFF64E;
		10'h5C: dout <= #1 24'hFFF66C;
		10'h5D: dout <= #1 24'hFFF7C4;
		10'h5E: dout <= #1 24'hFFFDE5;
		10'h5F: dout <= #1 24'hFFFB37;
		10'h60: dout <= #1 24'hB52;
		10'h61: dout <= #1 24'h17A;
		10'h62: dout <= #1 24'h4A8;
		10'h63: dout <= #1 24'hFFF6F6;
		10'h64: dout <= #1 24'hFFF820;
		10'h65: dout <= #1 24'hDCF;
		10'h66: dout <= #1 24'hFFFEA0;
		10'h67: dout <= #1 24'h396;
		10'h68: dout <= #1 24'hEE7;
		10'h69: dout <= #1 24'h479;
		10'h6A: dout <= #1 24'hC44;
		10'h6B: dout <= #1 24'hFFFC11;
		10'h6C: dout <= #1 24'hFFF833;
		10'h6D: dout <= #1 24'hB4A;
		10'h6E: dout <= #1 24'hFFF18D;
		10'h6F: dout <= #1 24'hC0F;
		10'h70: dout <= #1 24'hFFF309;
		10'h71: dout <= #1 24'hFFF32B;
		10'h72: dout <= #1 24'hFFFEDA;
		10'h73: dout <= #1 24'h425;
		10'h74: dout <= #1 24'hFFEE46;
		10'h75: dout <= #1 24'hF7;
		10'h76: dout <= #1 24'hFFFDCD;
		10'h77: dout <= #1 24'hD1D;
		10'h78: dout <= #1 24'hFFFACC;
		10'h79: dout <= #1 24'h629;
		10'h7A: dout <= #1 24'h718;
		10'h7B: dout <= #1 24'hFFF478;
		10'h7C: dout <= #1 24'hFFFE7B;
		10'h7D: dout <= #1 24'hA02;
		10'h7E: dout <= #1 24'h40D;
		10'h7F: dout <= #1 24'hFFFD45;
		10'h80: dout <= #1 24'h4D6;
		10'h81: dout <= #1 24'h652;
		10'h82: dout <= #1 24'hFFF262;
		10'h83: dout <= #1 24'hFFF1AE;
		10'h84: dout <= #1 24'hFFEF48;
		10'h85: dout <= #1 24'hA91;
		10'h86: dout <= #1 24'hFFFF8F;
		10'h87: dout <= #1 24'hFFFDA9;
		10'h88: dout <= #1 24'h1D6;
		10'h89: dout <= #1 24'h28A;
		10'h8A: dout <= #1 24'h5C4;
		10'h8B: dout <= #1 24'h10A9;
		10'h8C: dout <= #1 24'hBF4;
		10'h8D: dout <= #1 24'hC1B;
		10'h8E: dout <= #1 24'hFFFF09;
		10'h8F: dout <= #1 24'h227;
		10'h90: dout <= #1 24'h370;
		10'h91: dout <= #1 24'hFFFC5B;
		10'h92: dout <= #1 24'hFFFB54;
		10'h93: dout <= #1 24'h4DE;
		10'h94: dout <= #1 24'hFFFD16;
		10'h95: dout <= #1 24'hFFFFA8;
		10'h96: dout <= #1 24'h93D;
		10'h97: dout <= #1 24'h4A8;
		10'h98: dout <= #1 24'hFFFED5;
		10'h99: dout <= #1 24'hFFFFE1;
		10'h9A: dout <= #1 24'hFFFC68;
		10'h9B: dout <= #1 24'hFFF3AB;
		10'h9C: dout <= #1 24'hFFFB30;
		10'h9D: dout <= #1 24'hFFFDBE;
		10'h9E: dout <= #1 24'hFFF445;
		10'h9F: dout <= #1 24'hFFF1B8;
		10'hA0: dout <= #1 24'h6C2;
		10'hA1: dout <= #1 24'hFFFCA0;
		10'hA2: dout <= #1 24'hFFFBAD;
		10'hA3: dout <= #1 24'hFFFF0C;
		10'hA4: dout <= #1 24'h39E;
		10'hA5: dout <= #1 24'h408;
		10'hA6: dout <= #1 24'h1EF;
		10'hA7: dout <= #1 24'hFFF86B;
		10'hA8: dout <= #1 24'h832;
		10'hA9: dout <= #1 24'h3E6;
		10'hAA: dout <= #1 24'hFFF6D1;
		10'hAB: dout <= #1 24'h437;
		10'hAC: dout <= #1 24'hFFFE3B;
		10'hAD: dout <= #1 24'hFFFB10;
		10'hAE: dout <= #1 24'hFFF609;
		10'hAF: dout <= #1 24'hFFF754;
		10'hB0: dout <= #1 24'h90;
		10'hB1: dout <= #1 24'hFFFA35;
		10'hB2: dout <= #1 24'h72C;
		10'hB3: dout <= #1 24'h51;
		10'hB4: dout <= #1 24'h88A;
		10'hB5: dout <= #1 24'h31F;
		10'hB6: dout <= #1 24'hFFFB91;
		10'hB7: dout <= #1 24'hFFFE8B;
		10'hB8: dout <= #1 24'hFFFE40;
		10'hB9: dout <= #1 24'h49D;
		10'hBA: dout <= #1 24'h1F6;
		10'hBB: dout <= #1 24'hFFF005;
		10'hBC: dout <= #1 24'h9F3;
		10'hBD: dout <= #1 24'h103;
		10'hBE: dout <= #1 24'hFFFE05;
		10'hBF: dout <= #1 24'h46C;
		10'hC0: dout <= #1 24'hFFF9FB;
		10'hC1: dout <= #1 24'h110;
		10'hC2: dout <= #1 24'h5DD;
		10'hC3: dout <= #1 24'hFFFE63;
		10'hC4: dout <= #1 24'h3A5;
		10'hC5: dout <= #1 24'hFFFEE8;
		10'hC6: dout <= #1 24'hFFFED8;
		10'hC7: dout <= #1 24'h10;
		10'hC8: dout <= #1 24'hFFFE81;
		10'hC9: dout <= #1 24'hFFFDDE;
		10'hCA: dout <= #1 24'hFFF243;
		10'hCB: dout <= #1 24'hFFFC8E;
		10'hCC: dout <= #1 24'hFFFDF0;
		10'hCD: dout <= #1 24'hFFF4B2;
		10'hCE: dout <= #1 24'hFFFBF5;
		10'hCF: dout <= #1 24'h189;
		10'hD0: dout <= #1 24'h5D9;
		10'hD1: dout <= #1 24'h6B6;
		10'hD2: dout <= #1 24'h9;
		10'hD3: dout <= #1 24'h5C2;
		10'hD4: dout <= #1 24'hFFFE57;
		10'hD5: dout <= #1 24'h416;
		10'hD6: dout <= #1 24'hFFFC18;
		10'hD7: dout <= #1 24'h9C;
		10'hD8: dout <= #1 24'hFFF4D1;
		10'hD9: dout <= #1 24'h4FD;
		10'hDA: dout <= #1 24'hA03;
		10'hDB: dout <= #1 24'hFFF94A;
		10'hDC: dout <= #1 24'hFFFD9C;
		10'hDD: dout <= #1 24'h143;
		10'hDE: dout <= #1 24'hFFFE4D;
		10'hDF: dout <= #1 24'hFFF891;
		10'hE0: dout <= #1 24'h1A4;
		10'hE1: dout <= #1 24'hFFF49A;
		10'hE2: dout <= #1 24'hBAC;
		10'hE3: dout <= #1 24'hFFFE69;
		10'hE4: dout <= #1 24'h53B;
		10'hE5: dout <= #1 24'hFFFCAD;
		10'hE6: dout <= #1 24'h734;
		10'hE7: dout <= #1 24'hFFFFE7;
		10'hE8: dout <= #1 24'h308;
		10'hE9: dout <= #1 24'h4A2;
		10'hEA: dout <= #1 24'h4B7;
		10'hEB: dout <= #1 24'hFFF86F;
		10'hEC: dout <= #1 24'hFFF7DA;
		10'hED: dout <= #1 24'hFFFCA0;
		10'hEE: dout <= #1 24'h3FA;
		10'hEF: dout <= #1 24'hFFFCC6;
		10'hF0: dout <= #1 24'h2F4;
		10'hF1: dout <= #1 24'hFFFD65;
		10'hF2: dout <= #1 24'h662;
		10'hF3: dout <= #1 24'h1E7;
		10'hF4: dout <= #1 24'h4C0;
		10'hF5: dout <= #1 24'h18C;
		10'hF6: dout <= #1 24'h79;
		10'hF7: dout <= #1 24'h870;
		10'hF8: dout <= #1 24'hFFFED7;
		10'hF9: dout <= #1 24'h857;
		10'hFA: dout <= #1 24'h40A;
		10'hFB: dout <= #1 24'hFFF236;
		10'hFC: dout <= #1 24'hFFF5AB;
		10'hFD: dout <= #1 24'h2BF;
		10'hFE: dout <= #1 24'hFFF394;
		10'hFF: dout <= #1 24'hFFFB80;
		10'h100: dout <= #1 24'hFFE80E;
		10'h101: dout <= #1 24'hBA2;
		10'h102: dout <= #1 24'h1A5;
		10'h103: dout <= #1 24'h123;
		10'h104: dout <= #1 24'hFFF7B6;
		10'h105: dout <= #1 24'h3D8;
		10'h106: dout <= #1 24'h2E4;
		10'h107: dout <= #1 24'hFFFD01;
		10'h108: dout <= #1 24'hF9C;
		10'h109: dout <= #1 24'h680;
		10'h10A: dout <= #1 24'h456;
		10'h10B: dout <= #1 24'h25B;
		10'h10C: dout <= #1 24'h7E3;
		10'h10D: dout <= #1 24'h245;
		10'h10E: dout <= #1 24'hFFFF8B;
		10'h10F: dout <= #1 24'h1ED;
		10'h110: dout <= #1 24'hFFFE08;
		10'h111: dout <= #1 24'hFFFBD5;
		10'h112: dout <= #1 24'h507;
		10'h113: dout <= #1 24'h22C;
		10'h114: dout <= #1 24'hFFF22C;
		10'h115: dout <= #1 24'h94C;
		10'h116: dout <= #1 24'hFFF9B3;
		10'h117: dout <= #1 24'h37;
		10'h118: dout <= #1 24'hFFFA12;
		10'h119: dout <= #1 24'hFFF518;
		10'h11A: dout <= #1 24'hFFF752;
		10'h11B: dout <= #1 24'h62B;
		10'h11C: dout <= #1 24'hACE;
		10'h11D: dout <= #1 24'hFFF827;
		10'h11E: dout <= #1 24'hFFFBB5;
		10'h11F: dout <= #1 24'hFFF55B;
		10'h120: dout <= #1 24'hFFF26D;
		10'h121: dout <= #1 24'h18D;
		10'h122: dout <= #1 24'h9F;
		10'h123: dout <= #1 24'hFFFF02;
		10'h124: dout <= #1 24'h428;
		10'h125: dout <= #1 24'h250;
		10'h126: dout <= #1 24'h129;
		10'h127: dout <= #1 24'hFFFEA6;
		10'h128: dout <= #1 24'h75;
		10'h129: dout <= #1 24'h1767;
		10'h12A: dout <= #1 24'hFFF111;
		10'h12B: dout <= #1 24'hE56;
		10'h12C: dout <= #1 24'hFFFF8F;
		10'h12D: dout <= #1 24'hA24;
		10'h12E: dout <= #1 24'h3C7;
		10'h12F: dout <= #1 24'hFFF88B;
		10'h130: dout <= #1 24'hFFF67B;
		10'h131: dout <= #1 24'hFFF3B4;
		10'h132: dout <= #1 24'hFFFCB6;
		10'h133: dout <= #1 24'h6C3;
		10'h134: dout <= #1 24'h36;
		10'h135: dout <= #1 24'hFFFB50;
		10'h136: dout <= #1 24'h9E4;
		10'h137: dout <= #1 24'hB1D;
		10'h138: dout <= #1 24'hFFFAC7;
		10'h139: dout <= #1 24'hFFFBD0;
		10'h13A: dout <= #1 24'hFFF880;
		10'h13B: dout <= #1 24'h5C8;
		10'h13C: dout <= #1 24'hFFF6A8;
		10'h13D: dout <= #1 24'hFFFF5A;
		10'h13E: dout <= #1 24'hFFFDC5;
		10'h13F: dout <= #1 24'h59E;
		10'h140: dout <= #1 24'hFFF632;
		10'h141: dout <= #1 24'hFFF8AF;
		10'h142: dout <= #1 24'hFFFAF1;
		10'h143: dout <= #1 24'h546;
		10'h144: dout <= #1 24'hFFFEA1;
		10'h145: dout <= #1 24'h7AE;
		10'h146: dout <= #1 24'h69;
		10'h147: dout <= #1 24'hFFFF20;
		10'h148: dout <= #1 24'hA28;
		10'h149: dout <= #1 24'hFFFCB8;
		10'h14A: dout <= #1 24'hFFF6C4;
		10'h14B: dout <= #1 24'hFFFCAE;
		10'h14C: dout <= #1 24'hFFF979;
		10'h14D: dout <= #1 24'h564;
		10'h14E: dout <= #1 24'h1407;
		10'h14F: dout <= #1 24'hFFFB78;
		10'h150: dout <= #1 24'hFFFFF6;
		10'h151: dout <= #1 24'h176;
		10'h152: dout <= #1 24'hFFF757;
		10'h153: dout <= #1 24'h5A4;
		10'h154: dout <= #1 24'hFFF9CA;
		10'h155: dout <= #1 24'h177;
		10'h156: dout <= #1 24'hFFEF8B;
		10'h157: dout <= #1 24'hFFFC33;
		10'h158: dout <= #1 24'hACD;
		10'h159: dout <= #1 24'h76F;
		10'h15A: dout <= #1 24'hFFF65B;
		10'h15B: dout <= #1 24'hFFFB4F;
		10'h15C: dout <= #1 24'hFFF639;
		10'h15D: dout <= #1 24'hFFFA75;
		10'h15E: dout <= #1 24'hFFFC95;
		10'h15F: dout <= #1 24'hFFE519;
		10'h160: dout <= #1 24'hFFF8EF;
		10'h161: dout <= #1 24'hFFF6CA;
		10'h162: dout <= #1 24'hFFF6CD;
		10'h163: dout <= #1 24'h125D;
		10'h164: dout <= #1 24'hFFF64F;
		10'h165: dout <= #1 24'h4A1;
		10'h166: dout <= #1 24'hFFFDE7;
		10'h167: dout <= #1 24'hFFFD84;
		10'h168: dout <= #1 24'hFFF901;
		10'h169: dout <= #1 24'hFFF97B;
		10'h16A: dout <= #1 24'h44B;
		10'h16B: dout <= #1 24'h50C;
		10'h16C: dout <= #1 24'hFFFDC5;
		10'h16D: dout <= #1 24'hFFF686;
		10'h16E: dout <= #1 24'hFFFB00;
		10'h16F: dout <= #1 24'h37F;
		10'h170: dout <= #1 24'hFFFE38;
		10'h171: dout <= #1 24'hFFF767;
		10'h172: dout <= #1 24'h87A;
		10'h173: dout <= #1 24'h659;
		10'h174: dout <= #1 24'h3AA;
		10'h175: dout <= #1 24'h4B5;
		10'h176: dout <= #1 24'h5F3;
		10'h177: dout <= #1 24'hBCE;
		10'h178: dout <= #1 24'h87C;
		10'h179: dout <= #1 24'hFFF341;
		10'h17A: dout <= #1 24'hFFFF59;
		10'h17B: dout <= #1 24'h9EC;
		10'h17C: dout <= #1 24'h154;
		10'h17D: dout <= #1 24'h1F4;
		10'h17E: dout <= #1 24'hDC6;
		10'h17F: dout <= #1 24'h6C9;
		10'h180: dout <= #1 24'h82F;
		10'h181: dout <= #1 24'hFFF928;
		10'h182: dout <= #1 24'h15A;
		10'h183: dout <= #1 24'hFFF51E;
		10'h184: dout <= #1 24'h132;
		10'h185: dout <= #1 24'h127;
		10'h186: dout <= #1 24'h3F3;
		10'h187: dout <= #1 24'hFFF439;
		10'h188: dout <= #1 24'h676;
		10'h189: dout <= #1 24'hFFFE20;
		10'h18A: dout <= #1 24'h612;
		10'h18B: dout <= #1 24'hFFFC35;
		10'h18C: dout <= #1 24'h7FB;
		10'h18D: dout <= #1 24'hFFFDC3;
		10'h18E: dout <= #1 24'h996;
		10'h18F: dout <= #1 24'hFFF10C;
		10'h190: dout <= #1 24'hFFFC06;
		10'h191: dout <= #1 24'hFFFFC5;
		10'h192: dout <= #1 24'hFFFB42;
		10'h193: dout <= #1 24'hFFF56F;
		10'h194: dout <= #1 24'hFFF603;
		10'h195: dout <= #1 24'hFFF88E;
		10'h196: dout <= #1 24'hFFFDDB;
		10'h197: dout <= #1 24'h4EC;
		10'h198: dout <= #1 24'hFFF932;
		10'h199: dout <= #1 24'h3DF;
		10'h19A: dout <= #1 24'hFFEBCF;
		10'h19B: dout <= #1 24'hFFF952;
		10'h19C: dout <= #1 24'hFFF909;
		10'h19D: dout <= #1 24'h778;
		10'h19E: dout <= #1 24'h9C9;
		10'h19F: dout <= #1 24'hFFFDF4;
		10'h1A0: dout <= #1 24'hFFF519;
		10'h1A1: dout <= #1 24'hFFF732;
		10'h1A2: dout <= #1 24'hFFF4CB;
		10'h1A3: dout <= #1 24'h3F4;
		10'h1A4: dout <= #1 24'hFFF0C6;
		10'h1A5: dout <= #1 24'hFFFA77;
		10'h1A6: dout <= #1 24'h355;
		10'h1A7: dout <= #1 24'h150A;
		10'h1A8: dout <= #1 24'h631;
		10'h1A9: dout <= #1 24'h891;
		10'h1AA: dout <= #1 24'hF90;
		10'h1AB: dout <= #1 24'h359;
		10'h1AC: dout <= #1 24'hC93;
		10'h1AD: dout <= #1 24'hFFFFAF;
		10'h1AE: dout <= #1 24'hFFFD19;
		10'h1AF: dout <= #1 24'h3EE;
		10'h1B0: dout <= #1 24'hFFF883;
		10'h1B1: dout <= #1 24'h1F7;
		10'h1B2: dout <= #1 24'h76E;
		10'h1B3: dout <= #1 24'hFFFAAC;
		10'h1B4: dout <= #1 24'h285;
		10'h1B5: dout <= #1 24'h1DB;
		10'h1B6: dout <= #1 24'hFFF45B;
		10'h1B7: dout <= #1 24'h750;
		10'h1B8: dout <= #1 24'hFFF84C;
		10'h1B9: dout <= #1 24'h343;
		10'h1BA: dout <= #1 24'h5E4;
		10'h1BB: dout <= #1 24'h8F3;
		10'h1BC: dout <= #1 24'hFFFE04;
		10'h1BD: dout <= #1 24'h52A;
		10'h1BE: dout <= #1 24'h5E4;
		10'h1BF: dout <= #1 24'hFFFC38;
		10'h1C0: dout <= #1 24'h6EB;
		10'h1C1: dout <= #1 24'h4D7;
		10'h1C2: dout <= #1 24'h776;
		10'h1C3: dout <= #1 24'hFFFE72;
		10'h1C4: dout <= #1 24'h969;
		10'h1C5: dout <= #1 24'hFFFE5C;
		10'h1C6: dout <= #1 24'hF03;
		10'h1C7: dout <= #1 24'hFFFB9A;
		10'h1C8: dout <= #1 24'hFFFAA8;
		10'h1C9: dout <= #1 24'h557;
		10'h1CA: dout <= #1 24'hFFFBFD;
		10'h1CB: dout <= #1 24'hFFF00F;
		10'h1CC: dout <= #1 24'hC2C;
		10'h1CD: dout <= #1 24'hDCF;
		10'h1CE: dout <= #1 24'hFFF98F;
		10'h1CF: dout <= #1 24'h114B;
		10'h1D0: dout <= #1 24'hFFFF84;
		10'h1D1: dout <= #1 24'h2EC;
		10'h1D2: dout <= #1 24'hEF;
		10'h1D3: dout <= #1 24'h14D4;
		10'h1D4: dout <= #1 24'h348;
		10'h1D5: dout <= #1 24'hFFF997;
		10'h1D6: dout <= #1 24'hFFF0AC;
		10'h1D7: dout <= #1 24'h1001;
		10'h1D8: dout <= #1 24'h2C5;
		10'h1D9: dout <= #1 24'hFFF483;
		10'h1DA: dout <= #1 24'hFFF7B3;
		10'h1DB: dout <= #1 24'hFFF709;
		10'h1DC: dout <= #1 24'hFFFCFF;
		10'h1DD: dout <= #1 24'hFFF6D1;
		10'h1DE: dout <= #1 24'h97D;
		10'h1DF: dout <= #1 24'hFFFF39;
		10'h1E0: dout <= #1 24'hBA;
		10'h1E1: dout <= #1 24'h14DF;
		10'h1E2: dout <= #1 24'h809;
		10'h1E3: dout <= #1 24'h1D4;
		10'h1E4: dout <= #1 24'hD2;
		10'h1E5: dout <= #1 24'h91A;
		10'h1E6: dout <= #1 24'hFFF8F0;
		10'h1E7: dout <= #1 24'hFFF54B;
		10'h1E8: dout <= #1 24'h5BC;
		10'h1E9: dout <= #1 24'hFFFD2A;
		10'h1EA: dout <= #1 24'hDD6;
		10'h1EB: dout <= #1 24'hFFF6BF;
		10'h1EC: dout <= #1 24'hFFFCF4;
		10'h1ED: dout <= #1 24'hFFFD45;
		10'h1EE: dout <= #1 24'hFFF47C;
		10'h1EF: dout <= #1 24'h878;
		10'h1F0: dout <= #1 24'h49;
		10'h1F1: dout <= #1 24'hFFFB54;
		10'h1F2: dout <= #1 24'hFFF2E2;
		10'h1F3: dout <= #1 24'hFFF7D8;
		10'h1F4: dout <= #1 24'h32F;
		10'h1F5: dout <= #1 24'hFFFD40;
		10'h1F6: dout <= #1 24'h657;
		10'h1F7: dout <= #1 24'h366;
		10'h1F8: dout <= #1 24'h190B;
		10'h1F9: dout <= #1 24'hFFFCD3;
		10'h1FA: dout <= #1 24'h1ED;
		10'h1FB: dout <= #1 24'hFFFA30;
		10'h1FC: dout <= #1 24'h20A;
		10'h1FD: dout <= #1 24'hFFF8CA;
		10'h1FE: dout <= #1 24'hFFFE2E;
		10'h1FF: dout <= #1 24'hFDA;
		10'h200: dout <= #1 24'hBD4;
		10'h201: dout <= #1 24'h6F4;
		10'h202: dout <= #1 24'hFFF910;
		10'h203: dout <= #1 24'h203;
		10'h204: dout <= #1 24'h19F;
		10'h205: dout <= #1 24'h29B;
		10'h206: dout <= #1 24'h60F;
		10'h207: dout <= #1 24'h47D;
		10'h208: dout <= #1 24'hFFFF59;
		10'h209: dout <= #1 24'hFFFE5B;
		10'h20A: dout <= #1 24'h7F5;
		10'h20B: dout <= #1 24'h5E9;
		10'h20C: dout <= #1 24'hFFFD68;
		10'h20D: dout <= #1 24'hBF;
		10'h20E: dout <= #1 24'h3B0;
		10'h20F: dout <= #1 24'h167;
		10'h210: dout <= #1 24'hFFFC8D;
		10'h211: dout <= #1 24'h612;
		10'h212: dout <= #1 24'h8EF;
		10'h213: dout <= #1 24'hD5A;
		10'h214: dout <= #1 24'hA0F;
		10'h215: dout <= #1 24'h417;
		10'h216: dout <= #1 24'hFFFDDE;
		10'h217: dout <= #1 24'h5C8;
		10'h218: dout <= #1 24'h958;
		10'h219: dout <= #1 24'h132B;
		10'h21A: dout <= #1 24'hFFFE0A;
		10'h21B: dout <= #1 24'hE93;
		10'h21C: dout <= #1 24'hFFFB39;
		10'h21D: dout <= #1 24'hFFFFC4;
		10'h21E: dout <= #1 24'h787;
		10'h21F: dout <= #1 24'h3B2;
		10'h220: dout <= #1 24'h803;
		10'h221: dout <= #1 24'hFFFC0A;
		10'h222: dout <= #1 24'h506;
		10'h223: dout <= #1 24'h87A;
		10'h224: dout <= #1 24'h53C;
		10'h225: dout <= #1 24'hCE9;
		10'h226: dout <= #1 24'hFB5;
		10'h227: dout <= #1 24'hFFF038;
		10'h228: dout <= #1 24'hFFFDB6;
		10'h229: dout <= #1 24'hAF3;
		10'h22A: dout <= #1 24'h3B1;
		10'h22B: dout <= #1 24'h754;
		10'h22C: dout <= #1 24'hFFF892;
		10'h22D: dout <= #1 24'h197;
		10'h22E: dout <= #1 24'h3E9;
		10'h22F: dout <= #1 24'h1FD;
		10'h230: dout <= #1 24'h11F;
		10'h231: dout <= #1 24'hFFFA5A;
		10'h232: dout <= #1 24'h109A;
		10'h233: dout <= #1 24'hFE9;
		10'h234: dout <= #1 24'hC0E;
		10'h235: dout <= #1 24'hFFF76C;
		10'h236: dout <= #1 24'hFFFD91;
		10'h237: dout <= #1 24'h4CC;
		10'h238: dout <= #1 24'h5CB;
		10'h239: dout <= #1 24'hFFFB99;
		10'h23A: dout <= #1 24'h500;
		10'h23B: dout <= #1 24'h23C;
		10'h23C: dout <= #1 24'h29A;
		10'h23D: dout <= #1 24'hB46;
		10'h23E: dout <= #1 24'hFFFA57;
		10'h23F: dout <= #1 24'h772;
		10'h240: dout <= #1 24'h7D6;
		10'h241: dout <= #1 24'hB;
		10'h242: dout <= #1 24'h64B;
		10'h243: dout <= #1 24'h6D0;
		10'h244: dout <= #1 24'h1453;
		10'h245: dout <= #1 24'hFFFC45;
		10'h246: dout <= #1 24'hFFFEF5;
		10'h247: dout <= #1 24'hDF9;
		10'h248: dout <= #1 24'hAA2;
		10'h249: dout <= #1 24'h525;
		10'h24A: dout <= #1 24'h4D5;
		10'h24B: dout <= #1 24'h9F4;
		10'h24C: dout <= #1 24'hEF;
		10'h24D: dout <= #1 24'h247;
		10'h24E: dout <= #1 24'h27B;
		10'h24F: dout <= #1 24'h250;
		10'h250: dout <= #1 24'h841;
		10'h251: dout <= #1 24'hFFF8D1;
		10'h252: dout <= #1 24'hC97;
		10'h253: dout <= #1 24'h315;
		10'h254: dout <= #1 24'hFFFB57;
		10'h255: dout <= #1 24'hF5;
		10'h256: dout <= #1 24'hFFEFFE;
		10'h257: dout <= #1 24'hFFEFB5;
		10'h258: dout <= #1 24'h10B;
		10'h259: dout <= #1 24'hFFFB59;
		10'h25A: dout <= #1 24'h3EC;
		10'h25B: dout <= #1 24'hFFFBA5;
		10'h25C: dout <= #1 24'h4C7;
		10'h25D: dout <= #1 24'h95C;
		10'h25E: dout <= #1 24'hFFF933;
		10'h25F: dout <= #1 24'hFFFBE2;
		10'h260: dout <= #1 24'h3B3;
		10'h261: dout <= #1 24'h136;
		10'h262: dout <= #1 24'h64A;
		10'h263: dout <= #1 24'hAFD;
		10'h264: dout <= #1 24'hFFF0A5;
		10'h265: dout <= #1 24'h164;
		10'h266: dout <= #1 24'h232;
		10'h267: dout <= #1 24'hB4;
		10'h268: dout <= #1 24'hFFFDF7;
		10'h269: dout <= #1 24'hA26;
		10'h26A: dout <= #1 24'hFFF8AF;
		10'h26B: dout <= #1 24'hFFFDC1;
		10'h26C: dout <= #1 24'hFFF656;
		10'h26D: dout <= #1 24'hDDC;
		10'h26E: dout <= #1 24'hFFF7E2;
		10'h26F: dout <= #1 24'hFFF6FD;
		10'h270: dout <= #1 24'hFFFC47;
		10'h271: dout <= #1 24'h3F6;
		10'h272: dout <= #1 24'hFFFA27;
		10'h273: dout <= #1 24'h592;
		10'h274: dout <= #1 24'h11B3;
		10'h275: dout <= #1 24'h183;
		10'h276: dout <= #1 24'hFFFFF5;
		10'h277: dout <= #1 24'hFFF4E9;
		10'h278: dout <= #1 24'hFFFB79;
		10'h279: dout <= #1 24'hFFFD1F;
		10'h27A: dout <= #1 24'hFFF3AD;
		10'h27B: dout <= #1 24'h5BB;
		10'h27C: dout <= #1 24'h6AD;
		10'h27D: dout <= #1 24'hFFFF1C;
		10'h27E: dout <= #1 24'hFFF943;
		10'h27F: dout <= #1 24'hFFFD95;
		10'h280: dout <= #1 24'h400;
		10'h281: dout <= #1 24'hFFFE7A;
		10'h282: dout <= #1 24'hFFF41E;
		10'h283: dout <= #1 24'hFFFCB8;
		10'h284: dout <= #1 24'h89A;
		10'h285: dout <= #1 24'hBC5;
		10'h286: dout <= #1 24'hFFF09C;
		10'h287: dout <= #1 24'h3C6;
		10'h288: dout <= #1 24'h409;
		10'h289: dout <= #1 24'hFFFAAD;
		10'h28A: dout <= #1 24'hFFF4A2;
		10'h28B: dout <= #1 24'hFFF561;
		10'h28C: dout <= #1 24'hFFF365;
		10'h28D: dout <= #1 24'h9C;
		10'h28E: dout <= #1 24'h108;
		10'h28F: dout <= #1 24'h1513;
		10'h290: dout <= #1 24'hFFF8CC;
		10'h291: dout <= #1 24'hFFFCE6;
		10'h292: dout <= #1 24'h6A4;
		10'h293: dout <= #1 24'h113;
		10'h294: dout <= #1 24'hFFFEE0;
		10'h295: dout <= #1 24'h5B7;
		10'h296: dout <= #1 24'hFFF789;
		10'h297: dout <= #1 24'hFFFD7C;
		10'h298: dout <= #1 24'hFFFD5F;
		10'h299: dout <= #1 24'hFFF697;
		10'h29A: dout <= #1 24'h326;
		10'h29B: dout <= #1 24'hFFFE99;
		10'h29C: dout <= #1 24'h92E;
		10'h29D: dout <= #1 24'hFFF59E;
		10'h29E: dout <= #1 24'h7BF;
		10'h29F: dout <= #1 24'hFFFD97;
		10'h2A0: dout <= #1 24'hFFF8A8;
		10'h2A1: dout <= #1 24'hFFF6CE;
		10'h2A2: dout <= #1 24'h55B;
		10'h2A3: dout <= #1 24'h50C;
		10'h2A4: dout <= #1 24'hA89;
		10'h2A5: dout <= #1 24'hFFFB2C;
		10'h2A6: dout <= #1 24'hFFFC12;
		10'h2A7: dout <= #1 24'hFFF967;
		10'h2A8: dout <= #1 24'hFFF9BD;
		10'h2A9: dout <= #1 24'h84;
		10'h2AA: dout <= #1 24'h66;
		10'h2AB: dout <= #1 24'h77;
		10'h2AC: dout <= #1 24'h605;
		10'h2AD: dout <= #1 24'hFFFEE5;
		10'h2AE: dout <= #1 24'h161;
		10'h2AF: dout <= #1 24'h657;
		10'h2B0: dout <= #1 24'hFFFE08;
		10'h2B1: dout <= #1 24'hFFEC84;
		10'h2B2: dout <= #1 24'hBB;
		10'h2B3: dout <= #1 24'h200;
		10'h2B4: dout <= #1 24'h627;
		10'h2B5: dout <= #1 24'hBE7;
		10'h2B6: dout <= #1 24'hFFFEF8;
		10'h2B7: dout <= #1 24'h13D;
		10'h2B8: dout <= #1 24'hFFF1A0;
		10'h2B9: dout <= #1 24'hC14;
		10'h2BA: dout <= #1 24'hEB8;
		10'h2BB: dout <= #1 24'h289;
		10'h2BC: dout <= #1 24'h45A;
		10'h2BD: dout <= #1 24'hFFFC81;
		10'h2BE: dout <= #1 24'hFFF87D;
		10'h2BF: dout <= #1 24'hFFF267;
		10'h2C0: dout <= #1 24'h30;
		10'h2C1: dout <= #1 24'hFFF9F5;
		10'h2C2: dout <= #1 24'h133;
		10'h2C3: dout <= #1 24'hFFFA7E;
		10'h2C4: dout <= #1 24'hFFFF26;
		10'h2C5: dout <= #1 24'hFFFAFC;
		10'h2C6: dout <= #1 24'hFFFFE9;
		10'h2C7: dout <= #1 24'hFFFBBC;
		10'h2C8: dout <= #1 24'hFFF33D;
		10'h2C9: dout <= #1 24'hFFF89B;
		10'h2CA: dout <= #1 24'h3CF;
		10'h2CB: dout <= #1 24'h6;
		10'h2CC: dout <= #1 24'hFFFF04;
		10'h2CD: dout <= #1 24'hFFF8E3;
		10'h2CE: dout <= #1 24'hFFFFEE;
		10'h2CF: dout <= #1 24'h95F;
		10'h2D0: dout <= #1 24'h1AA;
		10'h2D1: dout <= #1 24'h2CF;
		10'h2D2: dout <= #1 24'hFFFC97;
		10'h2D3: dout <= #1 24'hFFF72F;
		10'h2D4: dout <= #1 24'h462;
		10'h2D5: dout <= #1 24'h649;
		10'h2D6: dout <= #1 24'hFFEF27;
		10'h2D7: dout <= #1 24'hFFFC51;
		10'h2D8: dout <= #1 24'hFFF073;
		10'h2D9: dout <= #1 24'hFFEE64;
		10'h2DA: dout <= #1 24'h754;
		10'h2DB: dout <= #1 24'hFFFAF6;
		10'h2DC: dout <= #1 24'hFFF6C0;
		10'h2DD: dout <= #1 24'h64C;
		10'h2DE: dout <= #1 24'h93D;
		10'h2DF: dout <= #1 24'h4BA;
		10'h2E0: dout <= #1 24'hB;
		10'h2E1: dout <= #1 24'h187;
		10'h2E2: dout <= #1 24'h3AE;
		10'h2E3: dout <= #1 24'hFFF84A;
		10'h2E4: dout <= #1 24'hB6D;
		10'h2E5: dout <= #1 24'hFFFB66;
		10'h2E6: dout <= #1 24'h4C4;
		10'h2E7: dout <= #1 24'hFFFD21;
		10'h2E8: dout <= #1 24'hAD6;
		10'h2E9: dout <= #1 24'hC24;
		10'h2EA: dout <= #1 24'hFFF45F;
		10'h2EB: dout <= #1 24'h709;
		10'h2EC: dout <= #1 24'h216;
		10'h2ED: dout <= #1 24'hFFF008;
		10'h2EE: dout <= #1 24'hFFF63F;
		10'h2EF: dout <= #1 24'hFFFC33;
		10'h2F0: dout <= #1 24'hFFF37C;
		10'h2F1: dout <= #1 24'hFFFA84;
		10'h2F2: dout <= #1 24'hFFFC91;
		10'h2F3: dout <= #1 24'hFFF733;
		10'h2F4: dout <= #1 24'hFFFC32;
		10'h2F5: dout <= #1 24'hD5;
		10'h2F6: dout <= #1 24'hFFFA0A;
		10'h2F7: dout <= #1 24'hFFFB4F;
		10'h2F8: dout <= #1 24'hFFF662;
		10'h2F9: dout <= #1 24'h292;
		10'h2FA: dout <= #1 24'hFFEB72;
		10'h2FB: dout <= #1 24'hFFF592;
		10'h2FC: dout <= #1 24'h9BB;
		10'h2FD: dout <= #1 24'hC77;
		10'h2FE: dout <= #1 24'hFFF776;
		10'h2FF: dout <= #1 24'hFFFA57;
		10'h300: dout <= #1 24'hFFFC3B;
		10'h301: dout <= #1 24'h5FF;
		10'h302: dout <= #1 24'hFFFB17;
		10'h303: dout <= #1 24'hFFEF08;
		10'h304: dout <= #1 24'h410;
		10'h305: dout <= #1 24'h93;
		10'h306: dout <= #1 24'h23C;
		10'h307: dout <= #1 24'h10C;
		10'h308: dout <= #1 24'hFFFB30;
		10'h309: dout <= #1 24'h130;
		10'h30A: dout <= #1 24'hFFF700;
		10'h30B: dout <= #1 24'h96D;
		10'h30C: dout <= #1 24'hFFFB6D;
		10'h30D: dout <= #1 24'h38;
		10'h30E: dout <= #1 24'hFFF656;
		10'h30F: dout <= #1 24'hFFF40A;
		10'h310: dout <= #1 24'h36C;
		10'h311: dout <= #1 24'h654;
		10'h312: dout <= #1 24'hFFF7F8;
		10'h313: dout <= #1 24'hFFF8F0;
		10'h314: dout <= #1 24'hFFFE0D;
		10'h315: dout <= #1 24'hFFFB2B;
		10'h316: dout <= #1 24'h5D9;
		10'h317: dout <= #1 24'hFFFD97;
		10'h318: dout <= #1 24'hFFF574;
		10'h319: dout <= #1 24'hFFFCAF;
		10'h31A: dout <= #1 24'hFFFFD2;
		10'h31B: dout <= #1 24'hFFF9BD;
		10'h31C: dout <= #1 24'h69F;
		10'h31D: dout <= #1 24'hFFFBEC;
		10'h31E: dout <= #1 24'hBA4;
		10'h31F: dout <= #1 24'hFFF4EA;
		10'h320: dout <= #1 24'hB6;
		10'h321: dout <= #1 24'h7A0;
		10'h322: dout <= #1 24'h38;
		10'h323: dout <= #1 24'h788;
		10'h324: dout <= #1 24'hFFF18E;
		10'h325: dout <= #1 24'h84E;
		10'h326: dout <= #1 24'hFFFAC2;
		10'h327: dout <= #1 24'h7F5;
		10'h328: dout <= #1 24'h2DF;
		10'h329: dout <= #1 24'h4A2;
		10'h32A: dout <= #1 24'hFFFDBE;
		10'h32B: dout <= #1 24'h380;
		10'h32C: dout <= #1 24'hFFFD81;
		10'h32D: dout <= #1 24'h139F;
		10'h32E: dout <= #1 24'h397;
		10'h32F: dout <= #1 24'hFFFDE4;
		10'h330: dout <= #1 24'hFFFE70;
		10'h331: dout <= #1 24'hFFF9C1;
		10'h332: dout <= #1 24'h8E2;
		10'h333: dout <= #1 24'hFFF7E5;
		10'h334: dout <= #1 24'hFFFAEB;
		10'h335: dout <= #1 24'h957;
		10'h336: dout <= #1 24'hA4D;
		10'h337: dout <= #1 24'h85;
		10'h338: dout <= #1 24'hFFF892;
		10'h339: dout <= #1 24'hE3;
		10'h33A: dout <= #1 24'hFFFAEC;
		10'h33B: dout <= #1 24'h495;
		10'h33C: dout <= #1 24'hFFF3EE;
		10'h33D: dout <= #1 24'h847;
		10'h33E: dout <= #1 24'h15B5;
		10'h33F: dout <= #1 24'h7A5;
		10'h340: dout <= #1 24'hFFFDE7;
		10'h341: dout <= #1 24'hFFF8E3;
		10'h342: dout <= #1 24'hFFFA75;
		10'h343: dout <= #1 24'hFFF6E4;
		10'h344: dout <= #1 24'hFFF450;
		10'h345: dout <= #1 24'h25;
		10'h346: dout <= #1 24'hFFEDA0;
		10'h347: dout <= #1 24'h7DC;
		10'h348: dout <= #1 24'hFFFFB9;
		10'h349: dout <= #1 24'hFFF826;
		10'h34A: dout <= #1 24'h5C7;
		10'h34B: dout <= #1 24'h714;
		10'h34C: dout <= #1 24'hFFFF2D;
		10'h34D: dout <= #1 24'h214;
		10'h34E: dout <= #1 24'hFFF542;
		10'h34F: dout <= #1 24'hFFFB1F;
		10'h350: dout <= #1 24'hFFF3D5;
		10'h351: dout <= #1 24'h254;
		10'h352: dout <= #1 24'hFFF86D;
		10'h353: dout <= #1 24'hFFF92C;
		10'h354: dout <= #1 24'hFFF7FA;
		10'h355: dout <= #1 24'hFFFEFA;
		10'h356: dout <= #1 24'h7AD;
		10'h357: dout <= #1 24'h2E7;
		10'h358: dout <= #1 24'h486;
		10'h359: dout <= #1 24'hFFFB80;
		10'h35A: dout <= #1 24'hFFFAE4;
		10'h35B: dout <= #1 24'hA1B;
		10'h35C: dout <= #1 24'hFEC;
		10'h35D: dout <= #1 24'hFFFFEB;
		10'h35E: dout <= #1 24'hFFF5D7;
		10'h35F: dout <= #1 24'hC2;
		10'h360: dout <= #1 24'hFFF89E;
		10'h361: dout <= #1 24'h574;
		10'h362: dout <= #1 24'hFFFAC1;
		10'h363: dout <= #1 24'hA5B;
		10'h364: dout <= #1 24'hA01;
		10'h365: dout <= #1 24'hB1C;
		10'h366: dout <= #1 24'hFFF5BD;
		10'h367: dout <= #1 24'hFFFC89;
		10'h368: dout <= #1 24'h13;
		10'h369: dout <= #1 24'hFFFB2C;
		10'h36A: dout <= #1 24'hFFFC13;
		10'h36B: dout <= #1 24'hFFF7E4;
		10'h36C: dout <= #1 24'h405;
		10'h36D: dout <= #1 24'hFFF3CA;
		10'h36E: dout <= #1 24'hFFF5EA;
		10'h36F: dout <= #1 24'h75A;
		10'h370: dout <= #1 24'h912;
		10'h371: dout <= #1 24'hFFF891;
		10'h372: dout <= #1 24'hFFFDFE;
		10'h373: dout <= #1 24'hFFFE3E;
		10'h374: dout <= #1 24'h231;
		10'h375: dout <= #1 24'hFFF79A;
		10'h376: dout <= #1 24'h60;
		10'h377: dout <= #1 24'hDCE;
		10'h378: dout <= #1 24'hFFF1B7;
		10'h379: dout <= #1 24'hFFF895;
		10'h37A: dout <= #1 24'h2C4;
		10'h37B: dout <= #1 24'h8A4;
		10'h37C: dout <= #1 24'hFFFA8E;
		10'h37D: dout <= #1 24'hFFF57B;
		10'h37E: dout <= #1 24'hFFF57D;
		10'h37F: dout <= #1 24'h305;
		10'h380: dout <= #1 24'hFFFD4B;
		10'h381: dout <= #1 24'hFFFF55;
		10'h382: dout <= #1 24'h48C;
		10'h383: dout <= #1 24'h8D2;
		10'h384: dout <= #1 24'hFFFF7C;
		10'h385: dout <= #1 24'hFFFAE3;
		10'h386: dout <= #1 24'h346;
		10'h387: dout <= #1 24'hFFF8EC;
		10'h388: dout <= #1 24'hFFF872;
		10'h389: dout <= #1 24'hC5B;
		10'h38A: dout <= #1 24'hFFFAB9;
		10'h38B: dout <= #1 24'h373;
		10'h38C: dout <= #1 24'h25F;
		10'h38D: dout <= #1 24'hFFF99C;
		10'h38E: dout <= #1 24'hFFFC92;
		10'h38F: dout <= #1 24'hFFFDAB;
		10'h390: dout <= #1 24'h317;
		10'h391: dout <= #1 24'hFFF23E;
		10'h392: dout <= #1 24'h71B;
		10'h393: dout <= #1 24'hFFFE55;
		10'h394: dout <= #1 24'h9F3;
		10'h395: dout <= #1 24'h412;
		10'h396: dout <= #1 24'h87D;
		10'h397: dout <= #1 24'hFFF43A;
		10'h398: dout <= #1 24'h66C;
		10'h399: dout <= #1 24'hFFF447;
		10'h39A: dout <= #1 24'h8B5;
		10'h39B: dout <= #1 24'hFFF7C3;
		10'h39C: dout <= #1 24'hE5F;
		10'h39D: dout <= #1 24'h102C;
		10'h39E: dout <= #1 24'hFFF573;
		10'h39F: dout <= #1 24'hFFF2FA;
		10'h3A0: dout <= #1 24'h755;
		10'h3A1: dout <= #1 24'hFFFE65;
		10'h3A2: dout <= #1 24'h5AC;
		10'h3A3: dout <= #1 24'h147A;
		10'h3A4: dout <= #1 24'h8D6;
		10'h3A5: dout <= #1 24'hFFFBE3;
		10'h3A6: dout <= #1 24'hFFF695;
		10'h3A7: dout <= #1 24'h19D;
		10'h3A8: dout <= #1 24'hFFF244;
		10'h3A9: dout <= #1 24'h837;
		10'h3AA: dout <= #1 24'h466;
		10'h3AB: dout <= #1 24'hFFFE29;
		10'h3AC: dout <= #1 24'hFFF5EE;
		10'h3AD: dout <= #1 24'h3AC;
		10'h3AE: dout <= #1 24'h232;
		10'h3AF: dout <= #1 24'h517;
		10'h3B0: dout <= #1 24'h83F;
		10'h3B1: dout <= #1 24'hFFFA33;
		10'h3B2: dout <= #1 24'hFFFA58;
		10'h3B3: dout <= #1 24'hFFF7C1;
		10'h3B4: dout <= #1 24'hFFFF2E;
		10'h3B5: dout <= #1 24'h7DE;
		10'h3B6: dout <= #1 24'hFFF47F;
		10'h3B7: dout <= #1 24'h29F;
		10'h3B8: dout <= #1 24'h375;
		10'h3B9: dout <= #1 24'hAC3;
		10'h3BA: dout <= #1 24'hFFF9C0;
		10'h3BB: dout <= #1 24'h96E;
		10'h3BC: dout <= #1 24'hFFFADF;
		10'h3BD: dout <= #1 24'h5F5;
		10'h3BE: dout <= #1 24'hFFF504;
		10'h3BF: dout <= #1 24'hFFF2DA;
		10'h3C0: dout <= #1 24'hFFF884;
		10'h3C1: dout <= #1 24'h76F;
		10'h3C2: dout <= #1 24'h11ED;
		10'h3C3: dout <= #1 24'hFFFD62;
		10'h3C4: dout <= #1 24'hFFF46B;
		10'h3C5: dout <= #1 24'hFFF71D;
		10'h3C6: dout <= #1 24'hE26;
		10'h3C7: dout <= #1 24'hFFF7C1;
		10'h3C8: dout <= #1 24'h706;
		10'h3C9: dout <= #1 24'hFFF072;
		10'h3CA: dout <= #1 24'h10F;
		10'h3CB: dout <= #1 24'hFFFEAA;
		10'h3CC: dout <= #1 24'hFFFD44;
		10'h3CD: dout <= #1 24'hADB;
		10'h3CE: dout <= #1 24'h4D9;
		10'h3CF: dout <= #1 24'hFFFDB9;
		10'h3D0: dout <= #1 24'hFFF5EC;
		10'h3D1: dout <= #1 24'h5F9;
		10'h3D2: dout <= #1 24'h124E;
		10'h3D3: dout <= #1 24'h9A9;
		10'h3D4: dout <= #1 24'hFFF623;
		10'h3D5: dout <= #1 24'h794;
		10'h3D6: dout <= #1 24'hFFF18D;
		10'h3D7: dout <= #1 24'h437;
		10'h3D8: dout <= #1 24'h5B0;
		10'h3D9: dout <= #1 24'h705;
		10'h3DA: dout <= #1 24'hA1;
		10'h3DB: dout <= #1 24'hFFFDE8;
		10'h3DC: dout <= #1 24'hFFFF9F;
		10'h3DD: dout <= #1 24'hFFF07F;
		10'h3DE: dout <= #1 24'hFFFFF9;
		10'h3DF: dout <= #1 24'h202;
		10'h3E0: dout <= #1 24'h32;
		10'h3E1: dout <= #1 24'hFFFECB;
		10'h3E2: dout <= #1 24'hA14;
		10'h3E3: dout <= #1 24'hFFFD67;
		10'h3E4: dout <= #1 24'h6E2;
		10'h3E5: dout <= #1 24'hA9;
		10'h3E6: dout <= #1 24'hFFF558;
		10'h3E7: dout <= #1 24'h8F6;
		10'h3E8: dout <= #1 24'hFFFEBF;
		10'h3E9: dout <= #1 24'hFFFDAA;
		10'h3EA: dout <= #1 24'hD96;
		10'h3EB: dout <= #1 24'h310;
		10'h3EC: dout <= #1 24'hBA5;
		10'h3ED: dout <= #1 24'hBB4;
		10'h3EE: dout <= #1 24'hFFF94A;
		10'h3EF: dout <= #1 24'hFFFF20;
		10'h3F0: dout <= #1 24'hFFFEE3;
		10'h3F1: dout <= #1 24'hFFF9B0;
		10'h3F2: dout <= #1 24'hFFFECB;
		10'h3F3: dout <= #1 24'hFFF621;
		10'h3F4: dout <= #1 24'hFFFB9B;
		10'h3F5: dout <= #1 24'hDFC;
		10'h3F6: dout <= #1 24'hFFF9F6;
		10'h3F7: dout <= #1 24'h7DB;
		10'h3F8: dout <= #1 24'h52;
		10'h3F9: dout <= #1 24'hD0E;
		10'h3FA: dout <= #1 24'h54A;
		10'h3FB: dout <= #1 24'h6AE;
		10'h3FC: dout <= #1 24'h390;
		10'h3FD: dout <= #1 24'h571;
		10'h3FE: dout <= #1 24'hFFFA68;
		10'h3FF: dout <= #1 24'h736;


    endcase

endmodule